/**74HC283 4?????? **/
module adder_4(
  input [3:0] A,         //??????
  input [3:0] B,         //??????
  input Cin,
  output [3:0] SUM,           //??????????????
  output Cout
);
  assign {Cout,SUM} = A + B +Cin;//????
endmodule
