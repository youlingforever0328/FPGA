module CD4532(input EI,input [7:0] I,output reg [2:0] Y,output reg GS,EO);
  integer k;
  always @(EI,I)
  begin
    if (EI == 0) begin Y = 3'd0; GS = 0;EO = 0;end
	else                 //?EI??1????????????
	   begin
	      GS = 1;EO = 0; //??????????????GS,EO????
		  for(k = 7;k >= 0;k = k - 1)
		    if(I[k]) begin Y = k; k = -1; end//???????????,k=-1??break??????????
		  if (I == 8'b00000000) begin Y = 3'd0;GS = 0;EO = 1; end//???????????
	   end 
  end
endmodule
